module CONTROL_INIT();
  task controlunit;
  // stuff
  endtask;
endmodule;
