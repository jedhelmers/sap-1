module ALU_INIT();
  task alu;
  // stuff
  endtask;
endmodule;
