module RAM_INIT();
  task ram;
  // stuff
  endtask;
endmodule;
