module OUT_7_SEGMENT_INIT();
  task 7_out;
  // stuff
  endtask;
endmodule;
