module REGISTER_INIT();
  task register;
  // stuff
  endtask;
endmodule;
