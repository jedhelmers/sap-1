module SAP1();
endmodule;
