module ram();
endmodule;
